`timescale 1ns / 1ps
// Full Adder
module FA(
output sum, cout, 
input a, b, cin
);
  wire w0, w1, w2;
  
  xor  (w0, a, b);
  xor  (sum, w0, cin);
  
  and  (w1, w0, cin);
  and  (w2, a, b);
  or  (cout, w1, w2);
endmodule
